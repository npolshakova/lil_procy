module add_four(four);

output [31:0] four;

assign four = 4;

endmodule